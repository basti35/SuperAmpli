** Profile: "SCHEMATIC1-V2_variabile"  [ X:\PROGETTO_ELETTRONICA\STADIO_2B\common_source-pspicefiles\schematic1\v2_variabile.sim ] 

** Creating circuit file "V2_variabile.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "X:\PROGETTO_ELETTRONICA\STADIO_2B\common_source-pspicefiles\schematic1\V2_variabile\V2_variabile_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.3_Demo\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 0.3ms 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
