** Profile: "SCHEMATIC1-time"  [ Y:\ORCAD\progetto\prove\stadio 3_caso a -pspicefiles\schematic1\time.sim ] 

** Creating circuit file "time.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../stadio 3_caso a -pspicefiles/pwrmos.lib" 
.LIB "../../../stadio 3_caso a -pspicefiles/stadio 3_caso a .lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.2\tools\PSpice\PSpice.ini file:

*Analysis directives: 
.TRAN  0 500us 0 1e-6 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
