** Profile: "SCHEMATIC1-Punto di lavoro"  [ Y:\ORCAD\PROGETTO\prove\stadio 3_caso a -PSpiceFiles\SCHEMATIC1\Punto di lavoro.sim ] 

** Creating circuit file "Punto di lavoro.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../stadio 3_caso a -pspicefiles/stadio 3_caso a .lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.2\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
