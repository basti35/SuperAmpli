** Profile: "SCHEMATIC1-tempo"  [ X:\PROGETTO_ELETTRONICA\STADIO_3\source_follower-pspicefiles\schematic1\tempo.sim ] 

** Creating circuit file "tempo.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.3_Demo\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10m 0 1u 
.OPTIONS STEPGMIN
.OPTIONS RELTOL= 1m
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
